module forwarding(input [2:0] rd_sw, input [2:0] lw_sw_sel, input [2:0] add_sel, input [2:0] sub_rm_sel,
	input [2:0] sub_rn_sel, input [2:0] cmp_shft_rd, input [2:0] EXMEM_rd1, input [2:0] MEMWB_rd1, input [2:0] MEMWB_rd2, 
	input EXMEM_regWrite1, input MEMWB_regWrite1, input MEMWB_regWrite2, input [1:0] ALUsrc1, input [1:0] ALUsrc2,
	input EXMEM_flagWrite1, input EXMEM_flagWrite2, input EXMEM_n_flag, output reg sel_n_flag, 
	output reg [1:0] sel_ALUsrc1, output reg [1:0] sel_ALUsrc2, output reg [1:0] sel_StoreData, output reg [1:0] sel_lw_sw_sel);
	
	//rs1 = storedatasel, lw_sw_sel = load/store address, add_sel = add, sub_rm_sel = sub, sub_rn_sel = sub/shift/cmp, cmp_shft_rd = shift/cmp
	//EXMEM_rd1 = write address of set1 instruction in ex/mem, rd12 = set2
	//MEMWB_rd1 = write address of set1 instruction in mem/wb, MEMWB_rd2 = set2
	//EXMEM_regWrite1 = regWrite of set1 instruction in ex/mem, regWrite12 = set2
	//MEMWB_regWrite1 = regWrite of set1 instruction in mem/wb, MEMWB_regWrite2 = set2
	//ALUsrc1 = aluALUsrc1 signal generated by ctrlckt, ALUsrc2 = aluALUsrc2
	
	always @(rd_sw or lw_sw_sel or add_sel or sub_rm_sel or sub_rn_sel or cmp_shft_rd or EXMEM_rd1 or MEMWB_rd1 or MEMWB_rd2 or ALUsrc1 or ALUsrc2 or EXMEM_flagWrite1 or EXMEM_flagWrite2 or EXMEM_regWrite1 or MEMWB_regWrite1 or MEMWB_regWrite2)
	begin
		sel_ALUsrc1 = 2'b00;
		sel_ALUsrc2 = 2'b00;
		//sel_EXMEMStoreData = 2'b00;
		sel_lw_sw_sel = 2'b00;
		sel_n_flag = 1'b0;
		sel_StoreData = 2'b00;
		
		if((EXMEM_regWrite1==1'b1) && (EXMEM_rd1==rd_sw)) sel_StoreData = 2'b01;
		else
		begin
		  // mem/wb1--store data dependency with g1
			if((MEMWB_regWrite1==1'b1) && (MEMWB_rd1==rd_sw)) sel_StoreData = 2'b10;			
     // mem/wb2--store data dependency with g2 load word
			if((MEMWB_regWrite2==1'b1) && (MEMWB_rd2==rd_sw)) sel_StoreData = 2'b11;
		end
		
		//address calculation dependency
		// ex/mem1--store/load address
		if((EXMEM_regWrite1==1'b1) && (EXMEM_rd1==lw_sw_sel)) sel_lw_sw_sel = 2'b01;
		else
		begin
		  // mem/wb1--store/load address dependency with g1
			if((MEMWB_regWrite1==1'b1) && (MEMWB_rd1==lw_sw_sel)) sel_lw_sw_sel = 2'b10;			
     // mem/wb2--store/load address dependency with g2 load word
			if((MEMWB_regWrite2==1'b1) && (MEMWB_rd2==lw_sw_sel)) sel_lw_sw_sel = 2'b11;
		end
		
		//ALU SRCA DEPENDENCY
		if((EXMEM_regWrite1==1'b1) && ((ALUsrc1==2'b00 && EXMEM_rd1==add_sel) || 
		   (ALUsrc1==2'b01 && EXMEM_rd1==sub_rn_sel) || 
		   (ALUsrc1==2'b10 && EXMEM_rd1==cmp_shft_rd))) sel_ALUsrc1 = 2'b01;// ex/mem1--aluALUsrc1
		else
		begin
			if((MEMWB_regWrite1==1'b1) && ((ALUsrc1==2'b00 && MEMWB_rd1==add_sel) || 
			   (ALUsrc1==2'b01 && MEMWB_rd1==sub_rn_sel) || 
			   (ALUsrc1==2'b10 && MEMWB_rd1==cmp_shft_rd))) sel_ALUsrc1 = 2'b10;// mem/wb1--aluALUsrc1
			
			if((MEMWB_regWrite2==1'b1) && ((ALUsrc1==2'b00 && MEMWB_rd2==add_sel) || 
			   (ALUsrc1==2'b01 && MEMWB_rd2==sub_rn_sel) || 
			   (ALUsrc1==2'b10 && MEMWB_rd2==cmp_shft_rd))) sel_ALUsrc1 = 2'b11;// mem/wb2--aluALUsrc1
		end
		
		//ALU SRCB DEPENDENCY.No condition check for add as it has only one source
		if((EXMEM_regWrite1==1'b1) && ((ALUsrc2==2'b00 && EXMEM_rd1==sub_rm_sel) ||
		   (ALUsrc2==2'b01 && EXMEM_rd1==sub_rn_sel))) sel_ALUsrc2 = 2'b01;// ex/mem1--aluALUsrc2
		else
		begin
			if((MEMWB_regWrite1==1'b1) && ((ALUsrc2==2'b00 && MEMWB_rd1==sub_rm_sel) || 
			  (ALUsrc2==2'b01 && MEMWB_rd1==sub_rn_sel))) sel_ALUsrc2 = 2'b10;// mem/wb1--aluALUsrc2
			
			if((MEMWB_regWrite2==1'b1) && ((ALUsrc2==2'b00 && MEMWB_rd2==sub_rm_sel) || 
			  (ALUsrc2==2'b01 && MEMWB_rd2==sub_rn_sel))) sel_ALUsrc2 = 2'b11;// mem/wb2--aluALUsrc2
		end
		
		/*??why EXMEM rdforlw_sw
		if((MEMWB_regWrite1==1'b1) && (MEMWB_rd1==EXMEM_rd_sw)) sel_EXMEMStoreData = 2'b01;// mem/wb aluOut
		if((MEMWB_regWrite2==1'b1) && (MEMWB_rd2==EXMEM_rd_sw)) sel_EXMEMStoreData = 2'b10;// mem/wb lw
		*/
		
		//flag forwarding.No need to frwd it from wb stage as we first write then read
		if((EXMEM_flagWrite1==1'b1) && ((EXMEM_n_flag==1'b1) || (EXMEM_flagWrite2==1'b0))) sel_n_flag = 1'b1; // EX/MEM
		
	end
endmodule

module forwarding_testbench;
  reg [2:0] EXMEM_rd_sw, lw_sw_sel, add_sel, sub_rm_sel, sub_rn_sel, cmp_shft_rd, EXMEM_rd1, MEMWB_rd1, MEMWB_rd2;
  reg EXMEM_regWrite1, MEMWB_regWrite1, MEMWB_regWrite2, EXMEM_n_flag;
  reg [1:0] ALUsrc1, ALUsrc2, EXMEM_flagWrite1,  EXMEM_flagWrite2;
  wire sel_n_flag, sel_ALUsrc1, sel_ALUsrc2, sel_EXMEMStoreData, sel_lw_sw_sel;
  forwarding forward(EXMEM_rd_sw, lw_sw_sel, add_sel, sub_rm_sel, sub_rn_sel, cmp_shft_rd, 
              EXMEM_rd1, MEMWB_rd1, MEMWB_rd2,EXMEM_regWrite1, MEMWB_regWrite1, MEMWB_regWrite2,
              ALUsrc1, ALUsrc2, EXMEM_flagWrite1, EXMEM_flagWrite2, sel_n_flag, sel_ALUsrc1, 
              sel_ALUsrc2, sel_EXMEMStoreData, sel_lw_sw_sel);
              
  
endmodule 